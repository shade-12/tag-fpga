
module tag_nios_system (
	bt_uart_RXD,
	bt_uart_TXD,
	clk_clk,
	hex_export,
	pll_locked_export,
	reset_reset_n,
	sd_card_b_SD_cmd,
	sd_card_b_SD_dat,
	sd_card_b_SD_dat3,
	sd_card_o_SD_clock,
	sdram_addr,
	sdram_ba,
	sdram_cas_n,
	sdram_cke,
	sdram_cs_n,
	sdram_dq,
	sdram_dqm,
	sdram_ras_n,
	sdram_we_n,
	sdram_clk_clk,
	wifi_uart_RXD,
	wifi_uart_TXD);	

	input		bt_uart_RXD;
	output		bt_uart_TXD;
	input		clk_clk;
	output	[6:0]	hex_export;
	output		pll_locked_export;
	input		reset_reset_n;
	inout		sd_card_b_SD_cmd;
	inout		sd_card_b_SD_dat;
	inout		sd_card_b_SD_dat3;
	output		sd_card_o_SD_clock;
	output	[12:0]	sdram_addr;
	output	[1:0]	sdram_ba;
	output		sdram_cas_n;
	output		sdram_cke;
	output		sdram_cs_n;
	inout	[15:0]	sdram_dq;
	output	[1:0]	sdram_dqm;
	output		sdram_ras_n;
	output		sdram_we_n;
	output		sdram_clk_clk;
	input		wifi_uart_RXD;
	output		wifi_uart_TXD;
endmodule
